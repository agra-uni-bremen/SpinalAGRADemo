module FirstModule
(
    input clk_i,
    input reset_i,
    input cond_i,
    output reg myRegister,
    output reg myRegisterWithReset
);

    wire 

endmodule
